module fetch();//stage 1

module execute();//stage 2

module generateparity();//stage 3

