`include "encoder.v"
`include "alu.v"
`include "parityGenerator.v"


module fetch(func,opcode);//stage 1
input [7:0] func;
output [2:0] opcode;
encoder


module execute();//stage 2

module generateparity();//stage 3

